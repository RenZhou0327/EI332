library verilog;
use verilog.vl_types.all;
entity sc_io_computer_vlg_vec_tst is
end sc_io_computer_vlg_vec_tst;
